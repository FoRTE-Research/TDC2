`timescale 1ns / 1ps

module my_not(
    input  a,
    output o
    );
    
    assign o = !a;

endmodule
