`timescale 1ns / 1ps

module my_and(
    input  a,
    input  b,
    output o
    );
    
    assign o = (a & b);

endmodule
